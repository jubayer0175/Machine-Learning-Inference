// platformniossdram.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module platformniossdram (
		input  wire        clk_clk,                           //          clk.clk
		output wire [31:0] hex_wire_export,                   //     hex_wire.export
		output wire [14:0] hps_0_ddr_mem_a,                   //    hps_0_ddr.mem_a
		output wire [2:0]  hps_0_ddr_mem_ba,                  //             .mem_ba
		output wire        hps_0_ddr_mem_ck,                  //             .mem_ck
		output wire        hps_0_ddr_mem_ck_n,                //             .mem_ck_n
		output wire        hps_0_ddr_mem_cke,                 //             .mem_cke
		output wire        hps_0_ddr_mem_cs_n,                //             .mem_cs_n
		output wire        hps_0_ddr_mem_ras_n,               //             .mem_ras_n
		output wire        hps_0_ddr_mem_cas_n,               //             .mem_cas_n
		output wire        hps_0_ddr_mem_we_n,                //             .mem_we_n
		output wire        hps_0_ddr_mem_reset_n,             //             .mem_reset_n
		inout  wire [31:0] hps_0_ddr_mem_dq,                  //             .mem_dq
		inout  wire [3:0]  hps_0_ddr_mem_dqs,                 //             .mem_dqs
		inout  wire [3:0]  hps_0_ddr_mem_dqs_n,               //             .mem_dqs_n
		output wire        hps_0_ddr_mem_odt,                 //             .mem_odt
		output wire [3:0]  hps_0_ddr_mem_dm,                  //             .mem_dm
		input  wire        hps_0_ddr_oct_rzqin,               //             .oct_rzqin
		output wire        hps_0_io_hps_io_emac1_inst_TX_CLK, //     hps_0_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_io_hps_io_emac1_inst_TXD0,   //             .hps_io_emac1_inst_TXD0
		output wire        hps_0_io_hps_io_emac1_inst_TXD1,   //             .hps_io_emac1_inst_TXD1
		output wire        hps_0_io_hps_io_emac1_inst_TXD2,   //             .hps_io_emac1_inst_TXD2
		output wire        hps_0_io_hps_io_emac1_inst_TXD3,   //             .hps_io_emac1_inst_TXD3
		input  wire        hps_0_io_hps_io_emac1_inst_RXD0,   //             .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_io_hps_io_emac1_inst_MDIO,   //             .hps_io_emac1_inst_MDIO
		output wire        hps_0_io_hps_io_emac1_inst_MDC,    //             .hps_io_emac1_inst_MDC
		input  wire        hps_0_io_hps_io_emac1_inst_RX_CTL, //             .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_io_hps_io_emac1_inst_TX_CTL, //             .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_io_hps_io_emac1_inst_RX_CLK, //             .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_io_hps_io_emac1_inst_RXD1,   //             .hps_io_emac1_inst_RXD1
		input  wire        hps_0_io_hps_io_emac1_inst_RXD2,   //             .hps_io_emac1_inst_RXD2
		input  wire        hps_0_io_hps_io_emac1_inst_RXD3,   //             .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_io_hps_io_qspi_inst_IO0,     //             .hps_io_qspi_inst_IO0
		inout  wire        hps_0_io_hps_io_qspi_inst_IO1,     //             .hps_io_qspi_inst_IO1
		inout  wire        hps_0_io_hps_io_qspi_inst_IO2,     //             .hps_io_qspi_inst_IO2
		inout  wire        hps_0_io_hps_io_qspi_inst_IO3,     //             .hps_io_qspi_inst_IO3
		output wire        hps_0_io_hps_io_qspi_inst_SS0,     //             .hps_io_qspi_inst_SS0
		output wire        hps_0_io_hps_io_qspi_inst_CLK,     //             .hps_io_qspi_inst_CLK
		inout  wire        hps_0_io_hps_io_sdio_inst_CMD,     //             .hps_io_sdio_inst_CMD
		inout  wire        hps_0_io_hps_io_sdio_inst_D0,      //             .hps_io_sdio_inst_D0
		inout  wire        hps_0_io_hps_io_sdio_inst_D1,      //             .hps_io_sdio_inst_D1
		output wire        hps_0_io_hps_io_sdio_inst_CLK,     //             .hps_io_sdio_inst_CLK
		inout  wire        hps_0_io_hps_io_sdio_inst_D2,      //             .hps_io_sdio_inst_D2
		inout  wire        hps_0_io_hps_io_sdio_inst_D3,      //             .hps_io_sdio_inst_D3
		inout  wire        hps_0_io_hps_io_usb1_inst_D0,      //             .hps_io_usb1_inst_D0
		inout  wire        hps_0_io_hps_io_usb1_inst_D1,      //             .hps_io_usb1_inst_D1
		inout  wire        hps_0_io_hps_io_usb1_inst_D2,      //             .hps_io_usb1_inst_D2
		inout  wire        hps_0_io_hps_io_usb1_inst_D3,      //             .hps_io_usb1_inst_D3
		inout  wire        hps_0_io_hps_io_usb1_inst_D4,      //             .hps_io_usb1_inst_D4
		inout  wire        hps_0_io_hps_io_usb1_inst_D5,      //             .hps_io_usb1_inst_D5
		inout  wire        hps_0_io_hps_io_usb1_inst_D6,      //             .hps_io_usb1_inst_D6
		inout  wire        hps_0_io_hps_io_usb1_inst_D7,      //             .hps_io_usb1_inst_D7
		input  wire        hps_0_io_hps_io_usb1_inst_CLK,     //             .hps_io_usb1_inst_CLK
		output wire        hps_0_io_hps_io_usb1_inst_STP,     //             .hps_io_usb1_inst_STP
		input  wire        hps_0_io_hps_io_usb1_inst_DIR,     //             .hps_io_usb1_inst_DIR
		input  wire        hps_0_io_hps_io_usb1_inst_NXT,     //             .hps_io_usb1_inst_NXT
		output wire        hps_0_io_hps_io_spim1_inst_CLK,    //             .hps_io_spim1_inst_CLK
		output wire        hps_0_io_hps_io_spim1_inst_MOSI,   //             .hps_io_spim1_inst_MOSI
		input  wire        hps_0_io_hps_io_spim1_inst_MISO,   //             .hps_io_spim1_inst_MISO
		output wire        hps_0_io_hps_io_spim1_inst_SS0,    //             .hps_io_spim1_inst_SS0
		input  wire        hps_0_io_hps_io_uart0_inst_RX,     //             .hps_io_uart0_inst_RX
		output wire        hps_0_io_hps_io_uart0_inst_TX,     //             .hps_io_uart0_inst_TX
		inout  wire        hps_0_io_hps_io_i2c0_inst_SDA,     //             .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_io_hps_io_i2c0_inst_SCL,     //             .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_io_hps_io_i2c1_inst_SDA,     //             .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_io_hps_io_i2c1_inst_SCL,     //             .hps_io_i2c1_inst_SCL
		input  wire [7:0]  key_wire_export,                   //     key_wire.export
		output wire [15:0] ledr_wire_export,                  //    ledr_wire.export
		output wire        pll_0_locked_export,               // pll_0_locked.export
		input  wire        reset_reset_n,                     //        reset.reset_n
		output wire        sdram_clk_clk,                     //    sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                   //   sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                     //             .ba
		output wire        sdram_wire_cas_n,                  //             .cas_n
		output wire        sdram_wire_cke,                    //             .cke
		output wire        sdram_wire_cs_n,                   //             .cs_n
		inout  wire [15:0] sdram_wire_dq,                     //             .dq
		output wire [1:0]  sdram_wire_dqm,                    //             .dqm
		output wire        sdram_wire_ras_n,                  //             .ras_n
		output wire        sdram_wire_we_n                    //             .we_n
	);

	wire         pll_0_outclk0_clk;                                           // pll_0:outclk_0 -> [irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, pio_0:clk, pio_1:clk, pio_2:clk, rst_controller:clk, timer_0:clk, timer_1:clk]
	wire         pll_0_outclk2_clk;                                           // pll_0:outclk_2 -> [mm_interconnect_0:pll_0_outclk2_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [26:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                  // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                                  // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                                 // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                                    // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                                 // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                  // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                                    // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                                 // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                 // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                 // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                 // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [31:0] hps_0_h2f_axi_master_wdata;                                  // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                                // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                                   // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                 // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                 // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                 // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                  // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                                // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [31:0] hps_0_h2f_axi_master_rdata;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                                // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                 // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                                 // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                                  // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                                   // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                                    // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                                 // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                 // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                                // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                                 // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect;                       // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                         // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                          // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                            // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                        // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_pio_1_s1_chipselect;                       // mm_interconnect_0:pio_1_s1_chipselect -> pio_1:chipselect
	wire  [31:0] mm_interconnect_0_pio_1_s1_readdata;                         // pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_1_s1_address;                          // mm_interconnect_0:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_0_pio_1_s1_write;                            // mm_interconnect_0:pio_1_s1_write -> pio_1:write_n
	wire  [31:0] mm_interconnect_0_pio_1_s1_writedata;                        // mm_interconnect_0:pio_1_s1_writedata -> pio_1:writedata
	wire  [31:0] mm_interconnect_0_pio_2_s1_readdata;                         // pio_2:readdata -> mm_interconnect_0:pio_2_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_2_s1_address;                          // mm_interconnect_0:pio_2_s1_address -> pio_2:address
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_1:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, pio_0:reset_n, pio_1:reset_n, pio_2:reset_n, rst_translator:in_reset, timer_0:reset_n, timer_1:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                                       // hps_0:h2f_rst_n -> rst_controller_002:reset_in0

	platformniossdram_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.h2f_mpu_eventi           (),                                  // h2f_mpu_events.eventi
		.h2f_mpu_evento           (),                                  //               .evento
		.h2f_mpu_standbywfe       (),                                  //               .standbywfe
		.h2f_mpu_standbywfi       (),                                  //               .standbywfi
		.mem_a                    (hps_0_ddr_mem_a),                   //         memory.mem_a
		.mem_ba                   (hps_0_ddr_mem_ba),                  //               .mem_ba
		.mem_ck                   (hps_0_ddr_mem_ck),                  //               .mem_ck
		.mem_ck_n                 (hps_0_ddr_mem_ck_n),                //               .mem_ck_n
		.mem_cke                  (hps_0_ddr_mem_cke),                 //               .mem_cke
		.mem_cs_n                 (hps_0_ddr_mem_cs_n),                //               .mem_cs_n
		.mem_ras_n                (hps_0_ddr_mem_ras_n),               //               .mem_ras_n
		.mem_cas_n                (hps_0_ddr_mem_cas_n),               //               .mem_cas_n
		.mem_we_n                 (hps_0_ddr_mem_we_n),                //               .mem_we_n
		.mem_reset_n              (hps_0_ddr_mem_reset_n),             //               .mem_reset_n
		.mem_dq                   (hps_0_ddr_mem_dq),                  //               .mem_dq
		.mem_dqs                  (hps_0_ddr_mem_dqs),                 //               .mem_dqs
		.mem_dqs_n                (hps_0_ddr_mem_dqs_n),               //               .mem_dqs_n
		.mem_odt                  (hps_0_ddr_mem_odt),                 //               .mem_odt
		.mem_dm                   (hps_0_ddr_mem_dm),                  //               .mem_dm
		.oct_rzqin                (hps_0_ddr_oct_rzqin),               //               .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_io_hps_io_emac1_inst_TX_CLK), //         hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_io_hps_io_emac1_inst_TXD0),   //               .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_io_hps_io_emac1_inst_TXD1),   //               .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_io_hps_io_emac1_inst_TXD2),   //               .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_io_hps_io_emac1_inst_TXD3),   //               .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_io_hps_io_emac1_inst_RXD0),   //               .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_io_hps_io_emac1_inst_MDIO),   //               .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_io_hps_io_emac1_inst_MDC),    //               .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_io_hps_io_emac1_inst_RX_CTL), //               .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_io_hps_io_emac1_inst_TX_CTL), //               .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_io_hps_io_emac1_inst_RX_CLK), //               .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_io_hps_io_emac1_inst_RXD1),   //               .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_io_hps_io_emac1_inst_RXD2),   //               .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_io_hps_io_emac1_inst_RXD3),   //               .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_io_hps_io_qspi_inst_IO0),     //               .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_io_hps_io_qspi_inst_IO1),     //               .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_io_hps_io_qspi_inst_IO2),     //               .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_io_hps_io_qspi_inst_IO3),     //               .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_io_hps_io_qspi_inst_SS0),     //               .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_io_hps_io_qspi_inst_CLK),     //               .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_io_hps_io_sdio_inst_CMD),     //               .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_io_hps_io_sdio_inst_D0),      //               .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_io_hps_io_sdio_inst_D1),      //               .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_io_hps_io_sdio_inst_CLK),     //               .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_io_hps_io_sdio_inst_D2),      //               .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_io_hps_io_sdio_inst_D3),      //               .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_io_hps_io_usb1_inst_D0),      //               .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_io_hps_io_usb1_inst_D1),      //               .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_io_hps_io_usb1_inst_D2),      //               .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_io_hps_io_usb1_inst_D3),      //               .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_io_hps_io_usb1_inst_D4),      //               .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_io_hps_io_usb1_inst_D5),      //               .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_io_hps_io_usb1_inst_D6),      //               .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_io_hps_io_usb1_inst_D7),      //               .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_io_hps_io_usb1_inst_CLK),     //               .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_io_hps_io_usb1_inst_STP),     //               .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_io_hps_io_usb1_inst_DIR),     //               .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_io_hps_io_usb1_inst_NXT),     //               .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_io_hps_io_spim1_inst_CLK),    //               .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_io_hps_io_spim1_inst_MOSI),   //               .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_io_hps_io_spim1_inst_MISO),   //               .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_io_hps_io_spim1_inst_SS0),    //               .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_io_hps_io_uart0_inst_RX),     //               .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_io_hps_io_uart0_inst_TX),     //               .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_io_hps_io_i2c0_inst_SDA),     //               .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_io_hps_io_i2c0_inst_SCL),     //               .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_io_hps_io_i2c1_inst_SDA),     //               .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_io_hps_io_i2c1_inst_SCL),     //               .hps_io_i2c1_inst_SCL
		.h2f_rst_n                (hps_0_h2f_reset_reset),             //      h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                           //  h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),         // h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),       //               .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),        //               .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),       //               .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),      //               .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),       //               .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),      //               .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),       //               .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),      //               .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),      //               .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),          //               .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),        //               .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),        //               .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),        //               .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),       //               .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),       //               .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),          //               .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),        //               .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),       //               .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),       //               .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),         //               .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),       //               .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),        //               .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),       //               .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),      //               .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),       //               .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),      //               .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),       //               .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),      //               .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),      //               .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),          //               .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),        //               .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),        //               .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),        //               .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),       //               .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready)        //               .rready
	);

	platformniossdram_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_0_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	platformniossdram_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_0_outclk0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	platformniossdram_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_0_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	platformniossdram_pio_0 pio_0 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (hex_wire_export)                        // external_connection.export
	);

	platformniossdram_pio_1 pio_1 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_1_s1_readdata),   //                    .readdata
		.out_port   (ledr_wire_export)                       // external_connection.export
	);

	platformniossdram_pio_2 pio_2 (
		.clk      (pll_0_outclk0_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_2_s1_readdata), //                    .readdata
		.in_port  (key_wire_export)                      // external_connection.export
	);

	platformniossdram_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),   // outclk0.clk
		.outclk_1 (sdram_clk_clk),       // outclk1.clk
		.outclk_2 (pll_0_outclk2_clk),   // outclk2.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	platformniossdram_sdram sdram (
		.clk            (pll_0_outclk2_clk),                        //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	platformniossdram_timer_0 timer_0 (
		.clk        (pll_0_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	platformniossdram_timer_0 timer_1 (
		.clk        (pll_0_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	platformniossdram_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                   //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                 //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                  //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                 //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                 //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                 //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                    //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                  //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                  //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                  //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                 //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                 //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                    //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                  //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                 //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                 //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                   //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                 //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                  //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                 //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                 //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                 //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                    //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                  //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                  //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                  //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                 //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                 //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                                     //                                                  clk_0_clk.clk
		.pll_0_outclk0_clk                                                (pll_0_outclk0_clk),                                           //                                              pll_0_outclk0.clk
		.pll_0_outclk2_clk                                                (pll_0_outclk2_clk),                                           //                                              pll_0_outclk2.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                              //                   nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset                          (rst_controller_001_reset_out_reset),                          //                          sdram_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                                 (nios2_gen2_0_data_master_address),                            //                                   nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                             (nios2_gen2_0_data_master_waitrequest),                        //                                                           .waitrequest
		.nios2_gen2_0_data_master_byteenable                              (nios2_gen2_0_data_master_byteenable),                         //                                                           .byteenable
		.nios2_gen2_0_data_master_read                                    (nios2_gen2_0_data_master_read),                               //                                                           .read
		.nios2_gen2_0_data_master_readdata                                (nios2_gen2_0_data_master_readdata),                           //                                                           .readdata
		.nios2_gen2_0_data_master_write                                   (nios2_gen2_0_data_master_write),                              //                                                           .write
		.nios2_gen2_0_data_master_writedata                               (nios2_gen2_0_data_master_writedata),                          //                                                           .writedata
		.nios2_gen2_0_data_master_debugaccess                             (nios2_gen2_0_data_master_debugaccess),                        //                                                           .debugaccess
		.nios2_gen2_0_instruction_master_address                          (nios2_gen2_0_instruction_master_address),                     //                            nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                      (nios2_gen2_0_instruction_master_waitrequest),                 //                                                           .waitrequest
		.nios2_gen2_0_instruction_master_read                             (nios2_gen2_0_instruction_master_read),                        //                                                           .read
		.nios2_gen2_0_instruction_master_readdata                         (nios2_gen2_0_instruction_master_readdata),                    //                                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                           .write
		.jtag_uart_0_avalon_jtag_slave_read                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                           .chipselect
		.nios2_gen2_0_debug_mem_slave_address                             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                               nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                                           .write
		.nios2_gen2_0_debug_mem_slave_read                                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                                           .read
		.nios2_gen2_0_debug_mem_slave_readdata                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                                           .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                                           .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                                           .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                                           .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                                           .debugaccess
		.onchip_memory2_0_s1_address                                      (mm_interconnect_0_onchip_memory2_0_s1_address),               //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                                           .clken
		.pio_0_s1_address                                                 (mm_interconnect_0_pio_0_s1_address),                          //                                                   pio_0_s1.address
		.pio_0_s1_write                                                   (mm_interconnect_0_pio_0_s1_write),                            //                                                           .write
		.pio_0_s1_readdata                                                (mm_interconnect_0_pio_0_s1_readdata),                         //                                                           .readdata
		.pio_0_s1_writedata                                               (mm_interconnect_0_pio_0_s1_writedata),                        //                                                           .writedata
		.pio_0_s1_chipselect                                              (mm_interconnect_0_pio_0_s1_chipselect),                       //                                                           .chipselect
		.pio_1_s1_address                                                 (mm_interconnect_0_pio_1_s1_address),                          //                                                   pio_1_s1.address
		.pio_1_s1_write                                                   (mm_interconnect_0_pio_1_s1_write),                            //                                                           .write
		.pio_1_s1_readdata                                                (mm_interconnect_0_pio_1_s1_readdata),                         //                                                           .readdata
		.pio_1_s1_writedata                                               (mm_interconnect_0_pio_1_s1_writedata),                        //                                                           .writedata
		.pio_1_s1_chipselect                                              (mm_interconnect_0_pio_1_s1_chipselect),                       //                                                           .chipselect
		.pio_2_s1_address                                                 (mm_interconnect_0_pio_2_s1_address),                          //                                                   pio_2_s1.address
		.pio_2_s1_readdata                                                (mm_interconnect_0_pio_2_s1_readdata),                         //                                                           .readdata
		.sdram_s1_address                                                 (mm_interconnect_0_sdram_s1_address),                          //                                                   sdram_s1.address
		.sdram_s1_write                                                   (mm_interconnect_0_sdram_s1_write),                            //                                                           .write
		.sdram_s1_read                                                    (mm_interconnect_0_sdram_s1_read),                             //                                                           .read
		.sdram_s1_readdata                                                (mm_interconnect_0_sdram_s1_readdata),                         //                                                           .readdata
		.sdram_s1_writedata                                               (mm_interconnect_0_sdram_s1_writedata),                        //                                                           .writedata
		.sdram_s1_byteenable                                              (mm_interconnect_0_sdram_s1_byteenable),                       //                                                           .byteenable
		.sdram_s1_readdatavalid                                           (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                                           .readdatavalid
		.sdram_s1_waitrequest                                             (mm_interconnect_0_sdram_s1_waitrequest),                      //                                                           .waitrequest
		.sdram_s1_chipselect                                              (mm_interconnect_0_sdram_s1_chipselect),                       //                                                           .chipselect
		.timer_0_s1_address                                               (mm_interconnect_0_timer_0_s1_address),                        //                                                 timer_0_s1.address
		.timer_0_s1_write                                                 (mm_interconnect_0_timer_0_s1_write),                          //                                                           .write
		.timer_0_s1_readdata                                              (mm_interconnect_0_timer_0_s1_readdata),                       //                                                           .readdata
		.timer_0_s1_writedata                                             (mm_interconnect_0_timer_0_s1_writedata),                      //                                                           .writedata
		.timer_0_s1_chipselect                                            (mm_interconnect_0_timer_0_s1_chipselect),                     //                                                           .chipselect
		.timer_1_s1_address                                               (mm_interconnect_0_timer_1_s1_address),                        //                                                 timer_1_s1.address
		.timer_1_s1_write                                                 (mm_interconnect_0_timer_1_s1_write),                          //                                                           .write
		.timer_1_s1_readdata                                              (mm_interconnect_0_timer_1_s1_readdata),                       //                                                           .readdata
		.timer_1_s1_writedata                                             (mm_interconnect_0_timer_1_s1_writedata),                      //                                                           .writedata
		.timer_1_s1_chipselect                                            (mm_interconnect_0_timer_1_s1_chipselect)                      //                                                           .chipselect
	);

	platformniossdram_irq_mapper irq_mapper (
		.clk           (pll_0_outclk0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk2_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
